// To Attatch to 0V Low 
module make_zero (w);
    output reg [15:0] w = 16'b0000;
endmodule
